module VirtualJTAG(input logic [1:0] ir_out,
                   input logic tdo,
                   output logic [1:0] ir_in,
                   output logic tck,
                   output logic tdi,
                   output logic virtual_state_cdr,
                   output logic virtual_state_cir,
                   output logic virtual_state_e1dr,
                   output logic virtual_state_e2dr,
                   output logic virtual_state_pdr,
                   output logic virtual_state_sdr,
                   output logic virtual_state_udr,
                   output logic virtual_state_uir);

sld_virtual_jtag	#(.sld_auto_instance_index("YES"),
                          .sld_instance_index(0),
                          .sld_ir_width(2),
                          .sld_sim_action(""),
                          .sld_sim_n_scan(0),
                          .sld_sim_total_length(0))
                        sld_virtual_jtag_component(.ir_out(ir_out),
                                                   .tdo(tdo),
                                                   .ir_in(ir_in),
                                                   .tck(tck),
                                                   .tdi(tdi),
                                                   .virtual_state_cdr(virtual_state_cdr),
                                                   .virtual_state_cir(virtual_state_cir),
                                                   .virtual_state_e1dr(virtual_state_e1dr),
                                                   .virtual_state_e2dr(virtual_state_e2dr),
                                                   .virtual_state_pdr(virtual_state_pdr),
                                                   .virtual_state_sdr(virtual_state_sdr),
                                                   .virtual_state_udr(virtual_state_udr),
                                                   .virtual_state_uir(virtual_state_uir),
                                                   .jtag_state_cdr(),
                                                   .jtag_state_cir(),
                                                   .jtag_state_e1dr(),
                                                   .jtag_state_e1ir(),
                                                   .jtag_state_e2dr(),
                                                   .jtag_state_e2ir(),
                                                   .jtag_state_pdr(),
                                                   .jtag_state_pir(),
                                                   .jtag_state_rti(),
                                                   .jtag_state_sdr(),
                                                   .jtag_state_sdrs(),
                                                   .jtag_state_sir(),
                                                   .jtag_state_sirs(),
                                                   .jtag_state_tlr(),
                                                   .jtag_state_udr(),
                                                   .jtag_state_uir(),
                                                   .tms());

endmodule
