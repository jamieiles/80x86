// Copyright Jamie Iles, 2017
//
// This file is part of s80x86.
//
// s80x86 is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
//
// s80x86 is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with s80x86.  If not, see <http://www.gnu.org/licenses/>.

module PosedgeToPulse(input logic clk,
                      input logic reset,
                      input logic d,
                      output logic q);

reg d_prev;

always_ff @(posedge clk)
    d_prev <= d;

always_ff @(posedge clk or posedge reset)
    if (reset) begin
        q <= 1'b0;
    end else begin
        q <= (d ^ d_prev) & d;
    end

endmodule
