`define CONFIG_SDRAM_SIZE (64 * 1024 * 1024)
`define CONFIG_VGA 1
`define CONFIG_PS2 1
`define CONFIG_NUM_LEDS 10
