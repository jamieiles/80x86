// Copyright Jamie Iles, 2017
//
// This file is part of s80x86.
//
// s80x86 is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
//
// s80x86 is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with s80x86.  If not, see <http://www.gnu.org/licenses/>.

`define CONFIG_SDRAM_SIZE (32 * 1024 * 1024)
`define CONFIG_VGA_DAC_BITS 4
`define CONFIG_VGA 1
`define CONFIG_PS2 1
`define CONFIG_NUM_LEDS 8
`define CONFIG_VIDEO_MEMORY_SIZE (16 * 1024)
`define CONFIG_SPEAKER 1
`define FORCE_M9K 1
