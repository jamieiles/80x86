`define CONFIG_SDRAM_SIZE (32 * 1024 * 1024)
`define CONFIG_LEDS
